package constants is

  -- Lattice iCEstick has a 12 Mhz oscillator
  constant clock_frequency : real := 12.0e6;

end package;

package body constants is

end package body;