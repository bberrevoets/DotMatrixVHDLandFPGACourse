library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity char_rom is
  port (
    clk : in std_logic;
    rst : in std_logic
  );
end char_rom;

architecture rtl of char_rom is

begin

end architecture;