library dot_matrix;
use dot_matrix.constants.all;

package sim_constants is

  constant clock_period : time := 1 sec / clock_frequency;

end package;
